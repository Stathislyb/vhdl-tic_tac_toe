library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity char_romx is
 port (
  address : in std_logic_vector(5 downto 0); 
  data : out std_logic_vector(63 downto 0));
end entity;

architecture RTLx of char_romx is
begin
  
 process(address)
 begin
  case address is
   when "000000" => data <= "1111100000000000000000000000000000000000000000000000000000011111";
   when "000001" => data <= "0111110000000000000000000000000000000000000000000000000000111110"; 
   when "000010" => data <= "0001111100000000000000000000000000000000000000000000000001111100"; 
   when "000011" => data <= "0000011111000000000000000000000000000000000000000000000001111100";
   when "000100" => data <= "0000000111110000000000000000000000000000000000000000000011111000"; 
   when "000101" => data <= "0000001111100000000000000000000000000000000000000000000111110000"; 
   when "000110" => data <= "0000000011111000000000000000000000000000000000000000001111100000"; 
   when "000111" => data <= "0000000000111110000000000000000000000000000000000000111110000000"; 
   when "001000" => data <= "0000000000011111000000000000000000000000000000000011111000000000"; 
   when "001001" => data <= "0000000000001111100000000000000000000000000000000111110000000000"; 
   when "001010" => data <= "0000000000000111110000000000000000000000000000000111110000000000"; 
   when "001011" => data <= "0000000000000001111100000000000000000000000000011111000000000000"; 
   when "001100" => data <= "0000000000000001111100000000000000000000000000111110000000000000"; 
   when "001101" => data <= "0000000000000000011111000000000000000000000011111000000000000000"; 
   when "001110" => data <= "0000000000000000001111100000000000000000000111110000000000000000"; 
   when "001111" => data <= "0000000000000000000111110000000000000000001111100000000000000000"; 
   when "010000" => data <= "0000000000000000000011111000000000000000011111000000000000000000"; 
   when "010001" => data <= "0000000000000000000001111100000000000001111100000000000000000000"; 
   when "010010" => data <= "0000000000000000000000111110000000000011111000000000000000000000"; 
   when "010011" => data <= "0000000000000000000000001111100000001111100000000000000000000000"; 
   when "010100" => data <= "0000000000000000000000000111110000011111000000000000000000000000"; 
   when "010101" => data <= "0000000000000000000000000011111001111100000000000000000000000000"; 
   when "010110" => data <= "0000000000000000000000000011111001111100000000000000000000000000"; 
   when "010111" => data <= "0000000000000000000000000000111111110000000000000000000000000000"; 
   when "011000" => data <= "0000000000000000000000000000001111100000000000000000000000000000"; 
   when "011001" => data <= "0000000000000000000000000000001111100000000000000000000000000000"; 
   when "011010" => data <= "0000000000000000000000000000111111100000000000000000000000000000"; 
   when "011011" => data <= "0000000000000000000000000001111101111000000000000000000000000000"; 
   when "011100" => data <= "0000000000000000000000000111110000111110000000000000000000000000"; 
   when "011101" => data <= "0000000000000000000000000111110000001111100000000000000000000000"; 
   when "011110" => data <= "0000000000000000000000011111000000001111100000000000000000000000"; 
   when "011111" => data <= "0000000000000000000000011111000000000011111000000000000000000000"; 
   when "100000" => data <= "0000000000000000000001111100000000000001111100000000000000000000"; 
   when "100001" => data <= "0000000000000000000001111100000000000000111110000000000000000000"; 
   when "100010" => data <= "0000000000000000000111110000000000000000001111100000000000000000"; 
   when "100011" => data <= "0000000000000000001111100000000000000000000011111000000000000000";
   when "100100" => data <= "0000000000000000011111000000000000000000000001111100000000000000"; 
   when "100101" => data <= "0000000000000001111100000000000000000000000000111110000000000000"; 
   when "100110" => data <= "0000000000000111110000000000000000000000000000001111100000000000"; 
   when "100111" => data <= "0000000000011111000000000000000000000000000000000111110000000000"; 
   when "101000" => data <= "0000000000111110000000000000000000000000000000000111110000000000"; 
   when "101001" => data <= "0000000011111000000000000000000000000000000000000001111100000000"; 
   when "101010" => data <= "0000000111110000000000000000000000000000000000000000111110000000"; 
   when "101011" => data <= "0000001111100000000000000000000000000000000000000000011111000000"; 
   when "101100" => data <= "0000011111000000000000000000000000000000000000000000001111100000"; 
   when "101101" => data <= "0001111100000000000000000000000000000000000000000000000011111000"; 
   when "101110" => data <= "0011111000000000000000000000000000000000000000000000000001111100"; 
   when "101111" => data <= "1111100000000000000000000000000000000000000000000000000000011111"; 
   when others => data <= "0000000000000000000000000000000000000000000000000000000000000000"; 
  end case;
 end process;

end RTLx;